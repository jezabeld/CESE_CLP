library IEEE;
use IEEE.std_logic_1164.all;

-- declaracion de entidad TEST BENCH
entity contNbmodMlento_tb is
end;

--cuerpo de arquitectura
architecture contNbmodMlento_tb_arq of contNbmodMlento_tb is
	-- seccion declarativa
	constant N_tb: natural := 5;
	constant M_tb: natural := 10;
	constant CICLOS_tb: natural :=4;

	signal clk_tb: std_logic := '0';
	signal rst_tb: std_logic := '1';
	signal ena_tb: std_logic := '1';
	signal q_tb: std_logic_vector (N_tb-1 downto 0);

begin
	-- seccion descriptiva
	clk_tb <= not clk_tb after 10 ns;
	rst_tb <= '0' after 25 ns;

	contNbmodMlento_inst: entity work.contNbmodMlento
		generic map(
			N => N_tb,
			M => M_tb,
			CICLOS => CICLOS_tb
		)
		port map(
			clk_i => clk_tb,
			rst_i => rst_tb,
			ena_i => ena_tb,
			q_o => q_tb 
		);
end;